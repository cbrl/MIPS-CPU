`ifndef ALU_OPS_SV
`define ALU_OPS_SV

typedef enum bit [3:0] {

	ALU_AND  = 4'b0000,
	ALU_OR   = 4'b0001,
	ALU_NOR  = 4'b0010,
	ALU_XOR  = 4'b0011,
	ALU_ADD  = 4'b0100,
	ALU_SUB  = 4'b0101,
	ALU_ADDU = 4'b0110,
	ALU_SUBU = 4'b0111,
	ALU_SLT  = 4'b1000,
	ALU_SLTU = 4'b1001,
	ALU_SGT  = 4'b1010,
	ALU_SGTU = 4'b1011,
	ALU_SLL  = 4'b1100,
	ALU_SRL  = 4'b1101,
	ALU_SRA  = 4'b1110,
	ALU_LUI  = 4'b1111

} ALU_OP;

`endif //ALU_OPS_SV
